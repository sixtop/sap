
module sap1 (
        //input wire clk,
        //input wire clr
    );

endmodule